library verilog;
use verilog.vl_types.all;
entity add_ress_sv_unit is
end add_ress_sv_unit;
