library verilog;
use verilog.vl_types.all;
entity nzp_comp_sv_unit is
end nzp_comp_sv_unit;
