library verilog;
use verilog.vl_types.all;
entity our_data_sv_unit is
end our_data_sv_unit;
