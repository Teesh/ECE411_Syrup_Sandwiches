library verilog;
use verilog.vl_types.all;
entity comp_tag_sv_unit is
end comp_tag_sv_unit;
