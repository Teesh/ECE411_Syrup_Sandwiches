library verilog;
use verilog.vl_types.all;
entity shift_ext_sv_unit is
end shift_ext_sv_unit;
