library verilog;
use verilog.vl_types.all;
entity add_ress is
    port(
        \in\            : in     vl_logic_vector(8 downto 0);
        index           : in     vl_logic_vector(2 downto 0);
        \out\           : out    vl_logic_vector(15 downto 0)
    );
end add_ress;
