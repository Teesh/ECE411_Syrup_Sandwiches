library verilog;
use verilog.vl_types.all;
entity masturgate_sv_unit is
end masturgate_sv_unit;
