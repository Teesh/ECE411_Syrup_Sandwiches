library verilog;
use verilog.vl_types.all;
entity ldb_shift_sv_unit is
end ldb_shift_sv_unit;
