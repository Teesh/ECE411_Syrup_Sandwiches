import lc3b_types::*;

module if_id
(
	input clk
);

register PC_reg
(
	.clk
);

register L_data
(
	.clk
);
endmodule: if_id
