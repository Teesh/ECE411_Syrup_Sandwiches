library verilog;
use verilog.vl_types.all;
entity mask2_sv_unit is
end mask2_sv_unit;
