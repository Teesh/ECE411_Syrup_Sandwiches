import lc3b_types::*;

module ldb_shift
(
	input clk,
	input logic [15:0] in,
	output logic [15:0] out
);


always_comb
begin


end
endmodule: ldb_shift