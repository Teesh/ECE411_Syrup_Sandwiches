module if_id
(

);