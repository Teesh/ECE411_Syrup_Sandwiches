library verilog;
use verilog.vl_types.all;
entity ryte_byte_sv_unit is
end ryte_byte_sv_unit;
