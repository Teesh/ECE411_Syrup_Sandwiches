import lc3b_types::*;

module shift_ext
(
	input clk,
	input logic [15:0] in,
	output logic [15:0] adj6_out, adj9_out, adj11_out, offset6_out, trapvect8_out, imm5_out, imm4_out
);

always_comb
begin

end
endmodule : shift_ext