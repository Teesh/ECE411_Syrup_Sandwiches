library verilog;
use verilog.vl_types.all;
entity br_enable_sv_unit is
end br_enable_sv_unit;
