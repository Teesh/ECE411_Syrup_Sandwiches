module if_id
(
	input clk
);

register PC_reg
(
	.clk
);