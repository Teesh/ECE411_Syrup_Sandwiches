library verilog;
use verilog.vl_types.all;
entity stb_shift_sv_unit is
end stb_shift_sv_unit;
